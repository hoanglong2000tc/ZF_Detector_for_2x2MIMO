module tb_ZF;
reg enable, clk, reset_n, accept_in;
wire accept_out, ready_out;

reg [255:0] H_matrix;
reg [127:0] y, n;
wire [127:0] X;

ZF uut(
    enable, clk, reset_n, accept_in, accept_out, ready_out, H_matrix, y, n, X
);

initial begin
    clk = 0;
    forever #5 clk = ~clk;
end
initial begin
    reset_n = 0; @(negedge clk);
    reset_n = 1;
end
initial begin
    enable = 1;
    accept_in = 1;
    #1950;
    enable = 0;
    #400;
    $stop;
end
reg [255:0] H_matrix_data[0:2];
initial begin
    
end

initial begin
    H_matrix_data[0] = 256'b0000101100110011000001001100110000001000000000001000100110011001100001001100110000001011001100110000100110011001000010000000000000000110011001101000101100110011000001100110011010001011001100110000101100110011000001100110011000001011001100110000011001100110;
    H_matrix_data[1] = 256'b0000111010111000100010110011001100001011001100111001100110011001000010110011001100001110101110000001100110011001000010110011001100000110011001101000111001100110000001100110011010001011001100110000111001100110000001100110011000001011001100110000011001100110;
    H_matrix_data[2] = 256'b0000011010111000100011001100110000001110011001101000100110011001000011001100110000000110101110000000100110011001000011100110011000001110011001101000110011001100000001100110011010001010000101000000110011001100000011100110011000001010000101000000011001100110;
end
initial begin
    y = 128'b00010000000000001000001100110011000000110011001100010000000000000000001100110011000001001100110010000100110011000000001100110011;
    n = 128'b00001000000000001000001001100110000000100110011000001000000000000001000000000000100100000000000000010000000000000001000000000000;
end
reg [1:0]i = 0;
always @(accept_out) begin
    if(accept_out) begin
        
        H_matrix = H_matrix_data[i];
        i = i + 1;
        if(i == 3) i = 0;
    end
end

endmodule

