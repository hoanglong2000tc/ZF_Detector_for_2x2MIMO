module tb_preprocess_ZF;
reg enable, clk, reset_n, accept_in;
wire accept_out, ready_out;
//
reg [127:0] y, n;
reg [255:0] invQ;
wire [127:0] Q_processed;

preprocess_ZF uut(enable, clk, reset_n, accept_in, accept_out, ready_out, y, n, invQ, Q_processed);

initial begin
    clk = 0;
    forever #5 clk = ~clk;
end
initial begin
    reset_n = 0; @(negedge clk);
    reset_n = 1;
end
initial begin
    enable = 1;
    accept_in = 1;
end

initial begin
    y = 128'b00010000000000001000001100110011000000110011001100010000000000000000001100110011000001001100110010000100110011000000001100110011;
    n = 128'b00001000000000001000001001100110000000100110011000001000000000000001000000000000100100000000000000010000000000000001000000000000;
end
reg [255:0] in [0 : 1];
initial begin
    in[0] = 256'b0000111010111000100010110011001100001011001100111001100110011001000010110011001100001110101110000001100110011001000010110011001100000110011001101000111001100110000001100110011010001011001100110000111001100110000001100110011000001011001100110000011001100110;
    in[1] = 256'b0001011010111000100011001100110000001110011001101000100110011001000011001100110000010110101110000000100110011001000011100110011000000110011001101000110011001100000001100110011010001010000101000000110011001100000001100110011000001010000101000000011001100110;
end
reg i = 0;
always @(accept_out) begin
    if(accept_out) begin
        invQ = in[i];
        i = i + 1;
    end
end



endmodule