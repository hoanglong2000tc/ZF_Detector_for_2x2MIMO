module transpose(
    output [255:0] out,
    input [255:0] in
);
assign out[255:240] = in[255:240];
assign out[239:224] = in[191:176];
assign out[191:176] = in[239:224];
assign out[223:208] = in[127:112];
assign out[127:112] = in[223:208];
assign out[207:192] = in[63:48];
assign out[63:48]   = in[207:192];
assign out[175:160] = in[175:160];
assign out[159:144] = in[111:96];
assign out[111:96]  = in[159:144];
assign out[143:128] = in[47:32];
assign out[47:32]   = in[143:128];
assign out[95:80] = in[95:80];
assign out[79:64]   = in[31:16];
assign out[31:16] = in[79:64];
assign out[15:0]    = in[15:0];

endmodule

// module tb_mul_4x4_4x2;
// reg clk, reset_n, start;
// wire done;
// wire [127:0]result;
// reg [255:0] A;
// reg[127:0] B;
// mul_4x4_4x2 uut(clk, reset_n, start, A, B, done, result);

// initial begin
//     clk = 0;
//     forever #5 clk = ~clk;
// end
// initial begin
//     reset_n = 0; @(negedge clk);
//     reset_n = 1;
// end
// initial begin
//     start = 0; repeat(2) @(negedge clk);
//     start = 1; @(negedge clk);
//     start = 0;
// end
// always @(done) begin
//     if(done) begin
//         repeat(5) @(negedge clk);
//         start = 1; @(negedge clk);
//         start = 0;
//     end
// end

// initial begin
//     A = 256'b0000001100110011100100000000000000001000000000001000100110011001000100000000000000000011001100110000100110011001000010000000000000000110011001101000101100110011000000011001100110000011001100110000101100110011000001100110011000000011001100110000000110011001;
//     B = 128'b00010000000000001000001100110011000000110011001100010000000000000000001100110011000001001100110010000100110011000000001100110011;
// end
// always @(result) begin
//     $display("%b",result);

// end
// endmodule
// //0000001100110011100100000000000000001000000000001000100110011001000100000000000000000011001100110000100110011001000010000000000000000110011001101000101100110011000000011001100110000011001100110000101100110011000001100110011000000011001100110000000110011001
// //100100000000000000001000000000001000100110011001000100000000000000000011001100110000100110011001000010000000000000000110011001101000101100110011000000011001100110000011001100110000101100110011000001100110011000000011001100110000000110011001