module tb_pipeline_QR_decomposition;
reg enable, clk, reset_n, accept_in;
wire accept_out, ready_out;

reg [511:0] H_matrix;
wire [511:0] Q_matrix, R_matrix;
QR uut(
    enable, clk, reset_n, accept_in, accept_out, ready_out, H_matrix, Q_matrix, R_matrix
);

initial begin
    clk = 0;
    forever #5 clk = ~clk;
end
initial begin
    reset_n = 0; @(negedge clk);
    reset_n = 1;
end
initial begin
    enable = 1;
    accept_in = 1;
end
reg [511:0] H_matrix_data[0:2];

initial begin
    H_matrix_data[0] = 512'b00000000101100110011001100110011000000000100110011001100110011010000000010000000000000000000000010000000100110011001100110011010100000000100110011001100110011010000000010110011001100110011001100000000100110011001100110011010000000001000000000000000000000000000000001100110011001100110011010000000101100110011001100110011000000000110011001100110011001101000000010110011001100110011001100000000101100110011001100110011000000000110011001100110011001100000000010110011001100110011001100000000011001100110011001100110;
    H_matrix_data[1] = 512'b00000000111010111000010100011111100000001011001100110011001100110000000010110011001100110011001110000001100110011001100110011010000000001011001100110011001100110000000011101011100001010001111100000001100110011001100110011010000000001011001100110011001100110000000001100110011001100110011010000000111001100110011001100110000000000110011001100110011001101000000010110011001100110011001100000000111001100110011001100110000000000110011001100110011001100000000010110011001100110011001100000000011001100110011001100110;
    H_matrix_data[2] = 512'b00000000011010111000010100011110100000001100110011001100110011010000000011100110011001100110011010000000100110011001100110011010000000001100110011001100110011010000000001101011100001010001111000000000100110011001100110011010000000001110011001100110011001100000000011100110011001100110011010000000110011001100110011001101000000000110011001100110011001101000000010100001010001111010111000000000110011001100110011001101000000001110011001100110011001100000000010100001010001111010111000000000011001100110011001100110;
end
reg [1:0]i = 0;
always @(accept_out) begin
    if(accept_out) begin
        
        H_matrix = H_matrix_data[i];
        i = i + 1;
        if(i == 3) i = 0;
    end
end

endmodule
